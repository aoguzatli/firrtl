module parameter_(
  input   always____,
  output  always$
);
  wire  assign__fork_;
  wire  edge__fork_;
  wire  always_ = ~always____;
  wire  always__ = always_;
  wire  always___ = 1'h0;
  endmodule__ assign_ (
    .fork_(assign__fork_)
  );
  endmodule_ edge_ (
    .fork_(edge__fork_)
  );
  assign always$ = 1'h0;
endmodule
module endmodule__(
  output  fork_
);
  wire [4:0] const_ = 5'h3;
  assign fork_ = 1'h1;
endmodule
module endmodule_(
  output  fork_
);
  wire [4:0] const_ = 5'h2;
  assign fork_ = 1'h0;
endmodule
