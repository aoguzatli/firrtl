// name:entries_info_ext depth:24 width:30 masked:false maskGran:30 maskSeg:1
module entries_info_ext(
  input R0_clk,
  input [4:0] R0_addr,
  input R0_en,
  output [29:0] R0_data,
  input W0_clk,
  input [4:0] W0_addr,
  input W0_en,
  input [29:0] W0_data
);



endmodule