// name:mem_ext depth:1024 width:16 masked:true maskGran:8 maskSeg:2
module mem_ext(
  input R0_clk,
  input [9:0] R0_addr,
  input R0_en,
  output [15:0] R0_data,
  input W0_clk,
  input [9:0] W0_addr,
  input W0_en,
  input [15:0] W0_data,
  input [1:0] W0_mask
);



endmodule