// name:mem_0_ext depth:7 width:16 masked:false maskGran:16 maskSeg:1
module mem_0_ext(
  input R0_clk,
  input [2:0] R0_addr,
  input R0_en,
  output [15:0] R0_data,
  input W0_clk,
  input [2:0] W0_addr,
  input W0_en,
  input [15:0] W0_data
);



endmodule