module Foo(
);
endmodule
